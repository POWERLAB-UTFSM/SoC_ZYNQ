module test (
    input aa,
    output wire bb,
);
    assign bb=aaa;
endmodule